ENTITY lshift_32_32 IS
PORT (
    D_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- Input 32-bit;
    D_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0) -- Output 32-bit;
  );
END lshift_32_32;
