ENTITY bus_merger IS
PORT (
    DATA_IN1 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    DATA_IN2 : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
    DATA_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END bus_merger;
